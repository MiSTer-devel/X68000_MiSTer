LIBRARY	IEEE;
USE	IEEE.STD_LOGIC_1164.ALL;
USE	IEEE.STD_LOGIC_UNSIGNED.ALL;

package FDC_sectinfo is

constant	nfmGap0		:integer	:=40;
constant	nmfmGap0	:integer	:=80;
constant	nfmSyncp	:integer	:=6;
constant	nmfmSyncp	:integer	:=12;
constant	nfmGap1		:integer	:=26;
constant	nmfmGap1	:integer	:=50;
constant	nfmSynci	:integer	:=6;
constant	nmfmSynci	:integer	:=12;
constant	nfmGap2		:integer	:=11;
constant	nmfmGap2	:integer	:=22;
constant	nfmSyncd	:integer	:=6;
constant	nmfmSyncd	:integer	:=12;

end FDC_sectinfo;

